../../src/verilog/opmem.sv