../../src/verilog/fp_add.sv