../../src/verilog/tb_fpu.sv