../../src/verilog/fpu.sv