module GraphPulse (
    input           clock,
    input           reset,
    input [15:0]    numVert,

    output          converge
);

endmodule // GraphPulse