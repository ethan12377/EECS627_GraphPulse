// TODO: implement PE in SV
