../../src/verilog/fp_div.sv