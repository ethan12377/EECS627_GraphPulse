../../src/verilog/fpuStim.sv