../../src/verilog/fp_mul.sv